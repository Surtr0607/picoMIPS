`define LIR 6'b000000
`define LSR 6'b000001
`define ADD 6'b000010
`define ADDI 6'b000011
`define MUL 6'b000100
`define MULI 6'b000101
`define WAIT0 6'b000110
`define WAIT1 6'b000111