//-----------------------------------------------------
// File Name   : alucodes.sv
// Function    : ALU module for picoMIPS
// Author:  Qi Zhong
// Last rev. 12 Mar 23
//-----------------------------------------------------


`define RA 2'b00
`define RB 2'b01
`define RADD 2'b10
`define RMUL 2'b11
